library verilog;
use verilog.vl_types.all;
entity Exercicio_Elevador is
    port(
        A               : in     vl_logic;
        B               : in     vl_logic;
        C               : in     vl_logic;
        D               : in     vl_logic;
        X               : out    vl_logic
    );
end Exercicio_Elevador;
