library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity flipflopd is
port
(

);

end entity;

architecture build of flipflopd is
begin




end architecture;