library verilog;
use verilog.vl_types.all;
entity Exercicio_Elevador_vlg_vec_tst is
end Exercicio_Elevador_vlg_vec_tst;
