library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity Exercicio_Elevador is
port
(
A, B, C, D : in std_logic;
X : out std_logic
);
end entity;

architecture build of Exercicio_Elevador is
begin
X <= (not A)AND(B OR D OR C);
end architecture;